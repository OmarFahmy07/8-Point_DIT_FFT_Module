// File : multiply.v
// Author : Omar Fahmy
// Date : 2/11/2022
// Version : 1
// Abstract : this file contains a fixed-point multiplication unit

//////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////// Module ports list, declaration, and data type ///////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////

module multiply #(parameter INT_WIDTH = 8,               // Integer Field Width
                  FRACT_WIDTH = 8,                       // Fractional Field Width
                  DATA_WIDTH = INT_WIDTH + FRACT_WIDTH)
                 (input wire [DATA_WIDTH-1 : 0] operand1,
                  input wire [DATA_WIDTH-1 : 0] operand2,
                  output reg [DATA_WIDTH-1 : 0] result);
    
    //////////////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////// Signals and Internal Connections ///////////////////////////////////
    //////////////////////////////////////////////////////////////////////////////////////////////////////
    
    reg [DATA_WIDTH-1 : 0] operand1_pos, operand2_pos;
    reg [2*DATA_WIDTH-1 : 0] mul_pos, mul;

    //////////////////////////////////////////////////////////////////////////////////////////////////////
    /////////////////////////////////////////// Procedural Blocks ////////////////////////////////////////
    //////////////////////////////////////////////////////////////////////////////////////////////////////
    
    always@(*)
    begin
        operand1_pos = operand1[DATA_WIDTH - 1] ? -operand1 : operand1;
        operand2_pos = operand2[DATA_WIDTH - 1] ? -operand2 : operand2;
        mul_pos      = operand1_pos * operand2_pos;
        mul          = operand1[DATA_WIDTH - 1] ^ operand2[DATA_WIDTH - 1] ? -mul_pos : mul_pos;
        result       = mul >> FRACT_WIDTH;
    end
    
endmodule
